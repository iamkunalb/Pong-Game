-- Bouncing Ball Video 
--
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;
USE  IEEE.STD_LOGIC_ARITH.all;
USE  IEEE.STD_LOGIC_UNSIGNED.all;
LIBRARY lpm;
USE lpm.lpm_components.ALL;

LIBRARY work;
USE work.de0core.all;

ENTITY bar IS
Generic(ADDR_WIDTH: integer := 12; DATA_WIDTH: integer := 1);

   PORT(SIGNAL PB1, PB2, Clock 			: IN std_logic;
        SIGNAL Red,Green,Blue 			: OUT std_logic;
        SIGNAL Horiz_sync,Vert_sync		: OUT std_logic);		
END bar;

architecture behavior of bar is

			-- Video Display Signals   
SIGNAL Red_Data, Green_Data, Blue_Data, vert_sync_int,
		reset, Ball_on, Direction			: std_logic;
SIGNAL Size 								: std_logic_vector(9 DOWNTO 0);  
SIGNAL Ball_Y_motion, Ball_X_motion : std_logic_vector(9 DOWNTO 0);
SIGNAL Ball_Y_pos, Ball_X_pos				: std_logic_vector(9 DOWNTO 0);
SIGNAL pixel_row, pixel_column				: std_logic_vector(9 DOWNTO 0); 

BEGIN           
   SYNC: vga_sync
 		PORT MAP(clock_25Mhz => clock, 
				red => red_data, green => green_data, blue => blue_data,	
    	     	red_out => red, green_out => green, blue_out => blue,
			 	horiz_sync_out => horiz_sync, vert_sync_out => vert_sync_int,
			 	pixel_row => pixel_row, pixel_column => pixel_column);

Size <= CONV_STD_LOGIC_VECTOR(8,10);
--Ball_X_pos <= CONV_STD_LOGIC_VECTOR(320,10);

		-- need internal copy of vert_sync to read
vert_sync <= vert_sync_int;

		-- Colors for pixel data on video signal
Red_Data <=  '1';
		-- Turn off Green and Blue when displaying ball
Green_Data <= NOT Ball_on;
Blue_Data <=  NOT Ball_on;

RGB_Display: Process (Ball_X_pos, Ball_Y_pos, pixel_column, pixel_row, Size)
BEGIN
			-- Set Ball_on ='1' to display ball
 IF ("00" & Ball_X_pos <= pixel_column + Size) AND
 			-- compare positive numbers only
 	("00" & Ball_X_pos + Size >= '0' & pixel_column) AND
	
 	('0' & Ball_Y_pos <= pixel_row + Size) AND
	
 	('0' & Ball_Y_pos + Size >= '0' & pixel_row ) THEN
 		Ball_on <= '1';
 	ELSE
 		Ball_on <= '0';

END IF;
END process RGB_Display;

Move_Ball: process
BEGIN
			-- Move ball once every vertical sync
	WAIT UNTIL vert_sync_int'event and vert_sync_int = '1';
	
	
			-- Bounce off top or bottom of screen
			IF ('0' & Ball_Y_pos) >= CONV_STD_LOGIC_VECTOR(480,10) - Size THEN
				Ball_Y_motion <= - CONV_STD_LOGIC_VECTOR(5,10);
			ELSIF Ball_Y_pos <= Size THEN
				Ball_Y_motion <= CONV_STD_LOGIC_VECTOR(5,10);
			END IF;
			
			IF ("00" & Ball_X_pos) >= CONV_STD_LOGIC_VECTOR(640,11) - Size THEN
				Ball_X_motion <= - CONV_STD_LOGIC_VECTOR(5,10);
			ELSIF("00" & Ball_X_pos) <= Size THEN
				Ball_X_motion <= CONV_STD_LOGIC_VECTOR(5,10);
			END IF;
			-- Compute next ball Y position
				Ball_X_pos <= Ball_X_pos + Ball_X_motion;
			
			-- Compute next ball Y position
				Ball_Y_pos <= Ball_Y_pos + Ball_Y_motion;
END process Move_Ball;


--	process(refresh_tick,ball_l,ball_t,xv_reg,yv_reg)
--	begin
--		ball_l_next <=ball_l;
--		ball_t_next <=ball_t;
--		xv_next<=xv_reg;
--		yv_next<=yv_reg;
--		if refresh_tick = '1' then
--			if ball_t> 400 and ball_l > (bar_l -ball_u) and ball_l < (bar_l +120)  then --top bar'a değdiği zaman
--				yv_next<= -y_v ;
--			elsif ball_t< 35  then--The ball hits the wall
--				yv_next<= y_v;
--			end if;
--			if ball_l < 10 then --The ball hits the left side of the screen
--				xv_next<= x_v;
--				elsif ball_l> 600 then                
--				xv_next<= -x_v ; --The ball hits the right side of the screen
--			end if; 
--			ball_l_next <=ball_l +xv_reg;
--			ball_t_next <=ball_t+yv_reg;               
--		end if;
--	end process;

END behavior;

